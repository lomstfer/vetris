module constants

pub const game_width = 10
pub const game_height = 20
pub const game_start_step_interval = 1.0 / 2.0
pub const game_acceleration_magic_number = 0.05