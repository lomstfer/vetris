module tetris

import irishgreencitrus.raylibv as r

struct Unit {
mut:
	x int
	y int
	color r.Color
}